// ID
module Sign_Extend(
    data_i,
    data_o
    );
               
// TO DO

          
endmodule