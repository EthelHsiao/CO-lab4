// ID
module Adder(
    src1_i,
	src2_i,
	sum_o
	);

// TO DO


endmodule                  